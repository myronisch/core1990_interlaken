-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- DO NOT EDIT THIS FILE
-- 
-- This file was generated from template '../firmware/sources/templates/pcie_package.vhd.template'
-- and register map registers-1.0.yaml, version 1.0
-- by the script 'wuppercodegen', version: 0.8.0,
-- using the following commandline:
-- 
-- ../software/wuppercodegen/wuppercodegen/cli.py registers-1.0.yaml ../firmware/sources/templates/pcie_package.vhd.template ../firmware/sources/packages/pcie_package.vhd
-- 
-- Please do NOT edit this file, but edit the source file at '../firmware/sources/templates/pcie_package.vhd.template'
-- 
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************
-- ***************************************************************************


--!------------------------------------------------------------------------------
--!
--!           NIKHEF - National Institute for Subatomic Physics
--!
--!                       Electronics Department
--!
--!-----------------------------------------------------------------------------
--! @class pcie_package
--!
--!
--! @author      Andrea Borga    (andrea.borga@nikhef.nl)<br>
--!              Frans Schreuder (frans.schreuder@nikhef.nl)
--!
--!
--! @date        07/01/2015    created
--!
--! @version     1.0
--!
--! @brief
--! This package contains the data types for the PCIe DMA core, as well as some
--! constants, addresses and register types for the application.
--!
--!
--! @detail
--!
--!-----------------------------------------------------------------------------
--! @TODO
--!
--!
--! ------------------------------------------------------------------------------
--! Virtex7 PCIe Gen3 DMA Core
--!
--! \copyright GNU LGPL License
--! Copyright (c) Nikhef, Amsterdam, All rights reserved. <br>
--! This library is free software; you can redistribute it and/or
--! modify it under the terms of the GNU Lesser General Public
--! License as published by the Free Software Foundation; either
--! version 3.0 of the License, or (at your option) any later version.
--! This library is distributed in the hope that it will be useful,
--! but WITHOUT ANY WARRANTY; without even the implied warranty of
--! MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the GNU
--! Lesser General Public License for more details.<br>
--! You should have received a copy of the GNU Lesser General Public
--! License along with this library.
--!

--! @brief ieee



library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_1164.all;

package pcie_package is

  function to_sl( A: std_logic_vector) return std_logic ;

  --
  -- PCIe DMA core: AXI-4 Stream interface
  type axis_type is record
    tdata   : std_logic_vector(255 downto 0);
    tkeep   : std_logic_vector(7 downto 0);
    tlast   : std_logic;
    tvalid  : std_logic;
  end record;

  type axis_r_type is record
    tready: std_logic;
  end record;

  --
  -- PCIe DMA core: descriptors
  type dma_descriptor_type is record
    start_address   : std_logic_vector(63 downto 0);
    current_address : std_logic_vector(63 downto 0);
    end_address     : std_logic_vector(63 downto 0);
    dword_count     : std_logic_vector(10 downto 0);
    read_not_write  : std_logic;     --1 means this is a read descriptor, 0: write descriptor
    enable          : std_logic;     --descriptor is valid
    wrap_around     : std_logic;     --1 means when end is reached, keep enabled and start over
    evencycle_dma   : std_logic;     --For every time the current_address overflows, this bit toggles
    evencycle_pc    : std_logic;     --For every time the pc pointer overflows, this bit toggles.
    pc_pointer      : std_logic_vector(63 downto 0); --Last address that the PC has read / written. For write: overflow and read until this cycle.
  end record;

  type dma_descriptors_type is array (natural range <>) of dma_descriptor_type;

  type dma_status_type is record
    descriptor_done: std_logic;  -- means the dma_descriptor in the array above has been handled, the enable field should then be cleared.
  end record;

  type dma_statuses_type is array(natural range <>) of dma_status_type;

  --
  -- PCIe DMA core: Interrupt Vectors
  type interrupt_vector_type is record
    int_vec_add  : std_logic_vector(63 downto 0);
    int_vec_data : std_logic_vector(31 downto 0);
    int_vec_ctrl : std_logic_vector(31 downto 0);
  end record;

  type interrupt_vectors_type is array (natural range <>) of interrupt_vector_type;

  --! Address Offset assignment
  --! --> BAR0 User Application Registers Addresses
  -- ### BAR0 registers: start
  constant REG_DESCRIPTOR_0        : std_logic_vector(19 downto 0) := x"00000";
  constant REG_DESCRIPTOR_0a       : std_logic_vector(19 downto 0) := x"00010";
  constant REG_DESCRIPTOR_1        : std_logic_vector(19 downto 0) := x"00020";
  constant REG_DESCRIPTOR_1a       : std_logic_vector(19 downto 0) := x"00030";
  constant REG_DESCRIPTOR_2        : std_logic_vector(19 downto 0) := x"00040";
  constant REG_DESCRIPTOR_2a       : std_logic_vector(19 downto 0) := x"00050";
  constant REG_DESCRIPTOR_3        : std_logic_vector(19 downto 0) := x"00060";
  constant REG_DESCRIPTOR_3a       : std_logic_vector(19 downto 0) := x"00070";
  constant REG_DESCRIPTOR_4        : std_logic_vector(19 downto 0) := x"00080";
  constant REG_DESCRIPTOR_4a       : std_logic_vector(19 downto 0) := x"00090";
  constant REG_DESCRIPTOR_5        : std_logic_vector(19 downto 0) := x"000A0";
  constant REG_DESCRIPTOR_5a       : std_logic_vector(19 downto 0) := x"000B0";
  constant REG_DESCRIPTOR_6        : std_logic_vector(19 downto 0) := x"000C0";
  constant REG_DESCRIPTOR_6a       : std_logic_vector(19 downto 0) := x"000D0";
  constant REG_DESCRIPTOR_7        : std_logic_vector(19 downto 0) := x"000E0";
  constant REG_DESCRIPTOR_7a       : std_logic_vector(19 downto 0) := x"000F0";
  constant REG_DESCRIPTOR_8        : std_logic_vector(19 downto 0) := x"00100";
  constant REG_DESCRIPTOR_8a       : std_logic_vector(19 downto 0) := x"00110";
  constant REG_DESCRIPTOR_9        : std_logic_vector(19 downto 0) := x"00120";
  constant REG_DESCRIPTOR_9a       : std_logic_vector(19 downto 0) := x"00130";
  constant REG_DESCRIPTOR_10       : std_logic_vector(19 downto 0) := x"00140";
  constant REG_DESCRIPTOR_10a      : std_logic_vector(19 downto 0) := x"00150";
  constant REG_DESCRIPTOR_11       : std_logic_vector(19 downto 0) := x"00160";
  constant REG_DESCRIPTOR_11a      : std_logic_vector(19 downto 0) := x"00170";
  constant REG_DESCRIPTOR_12       : std_logic_vector(19 downto 0) := x"00180";
  constant REG_DESCRIPTOR_12a      : std_logic_vector(19 downto 0) := x"00190";
  constant REG_DESCRIPTOR_13       : std_logic_vector(19 downto 0) := x"001A0";
  constant REG_DESCRIPTOR_13a      : std_logic_vector(19 downto 0) := x"001B0";
  constant REG_DESCRIPTOR_14       : std_logic_vector(19 downto 0) := x"001C0";
  constant REG_DESCRIPTOR_14a      : std_logic_vector(19 downto 0) := x"001D0";
  constant REG_DESCRIPTOR_15       : std_logic_vector(19 downto 0) := x"001E0";
  constant REG_DESCRIPTOR_15a      : std_logic_vector(19 downto 0) := x"001F0";
  constant REG_STATUS_0            : std_logic_vector(19 downto 0) := x"00200";
  constant REG_STATUS_1            : std_logic_vector(19 downto 0) := x"00210";
  constant REG_STATUS_2            : std_logic_vector(19 downto 0) := x"00220";
  constant REG_STATUS_3            : std_logic_vector(19 downto 0) := x"00230";
  constant REG_STATUS_4            : std_logic_vector(19 downto 0) := x"00240";
  constant REG_STATUS_5            : std_logic_vector(19 downto 0) := x"00250";
  constant REG_STATUS_6            : std_logic_vector(19 downto 0) := x"00260";
  constant REG_STATUS_7            : std_logic_vector(19 downto 0) := x"00270";
  constant REG_STATUS_8            : std_logic_vector(19 downto 0) := x"00280";
  constant REG_STATUS_9            : std_logic_vector(19 downto 0) := x"00290";
  constant REG_STATUS_10           : std_logic_vector(19 downto 0) := x"002A0";
  constant REG_STATUS_11           : std_logic_vector(19 downto 0) := x"002B0";
  constant REG_STATUS_12           : std_logic_vector(19 downto 0) := x"002C0";
  constant REG_STATUS_13           : std_logic_vector(19 downto 0) := x"002D0";
  constant REG_STATUS_14           : std_logic_vector(19 downto 0) := x"002E0";
  constant REG_STATUS_15           : std_logic_vector(19 downto 0) := x"002F0";
  constant REG_BAR0                : std_logic_vector(19 downto 0) := x"00300";
  constant REG_BAR1                : std_logic_vector(19 downto 0) := x"00310";
  constant REG_BAR2                : std_logic_vector(19 downto 0) := x"00320";
  constant REG_DESCRIPTOR_ENABLE   : std_logic_vector(19 downto 0) := x"00400";
  constant REG_FIFO_FLUSH          : std_logic_vector(19 downto 0) := x"00410";
  constant REG_DMA_RESET           : std_logic_vector(19 downto 0) := x"00420";
  constant REG_SOFT_RESET          : std_logic_vector(19 downto 0) := x"00430";
  constant REG_REGISTER_RESET      : std_logic_vector(19 downto 0) := x"00440";
  constant REG_FROMHOST_FULL_THRESH: std_logic_vector(19 downto 0) := x"00450";
  constant REG_TOHOST_FULL_THRESH  : std_logic_vector(19 downto 0) := x"00460";
  
  -- BAR0 registers: end

  --! Address Offset assignment
  --! --> BAR1 User Application Registers Addresses
  -- ### BAR1 registers: start
     -- interrupt vectors
  constant REG_INT_VEC_00          : std_logic_vector(19 downto 0) := x"00000";
  constant REG_INT_VEC_01          : std_logic_vector(19 downto 0) := x"00010";
  constant REG_INT_VEC_02          : std_logic_vector(19 downto 0) := x"00020";
  constant REG_INT_VEC_03          : std_logic_vector(19 downto 0) := x"00030";
  constant REG_INT_VEC_04          : std_logic_vector(19 downto 0) := x"00040";
  constant REG_INT_VEC_05          : std_logic_vector(19 downto 0) := x"00050";
  constant REG_INT_VEC_06          : std_logic_vector(19 downto 0) := x"00060";
  constant REG_INT_VEC_07          : std_logic_vector(19 downto 0) := x"00070";
  constant REG_INT_TAB_EN          : std_logic_vector(19 downto 0) := x"00100";
  -- BAR1 registers: end


  --! Address Offset assignment
  --! --> BAR2 User Application Registers Addresses
  --! -- leave 16x8 = 128 bits space per register
  ------------------------------------
  ---- ## GENERATED code BEGIN #1 ----
  ------------------------------------

  --** Bar2

  --** GenericBoardInformation
  constant REG_REG_MAP_VERSION                : std_logic_vector(19 downto 0) := x"00000";
  constant REG_BOARD_ID_TIMESTAMP             : std_logic_vector(19 downto 0) := x"00010";
  constant REG_BOARD_ID_SVN                   : std_logic_vector(19 downto 0) := x"00020";
  constant REG_STATUS_LEDS                    : std_logic_vector(19 downto 0) := x"00030";
  constant REG_GENERIC_CONSTANTS              : std_logic_vector(19 downto 0) := x"00040";
  constant REG_CARD_TYPE                      : std_logic_vector(19 downto 0) := x"00050";

  --** ApplicationSpecific
  constant REG_LFSR_SEED_0                    : std_logic_vector(19 downto 0) := x"01000";
  constant REG_LFSR_SEED_1                    : std_logic_vector(19 downto 0) := x"01010";
  constant REG_LFSR_SEED_2                    : std_logic_vector(19 downto 0) := x"01020";
  constant REG_LFSR_SEED_3                    : std_logic_vector(19 downto 0) := x"01030";
  constant REG_APP_MUX                        : std_logic_vector(19 downto 0) := x"01040";
  constant REG_LFSR_LOAD_SEED                 : std_logic_vector(19 downto 0) := x"01050";
  constant REG_APP_ENABLE                     : std_logic_vector(19 downto 0) := x"01060";

  --** HouseKeepingControlsAndMonitors
  constant REG_MMCM_MAIN_PLL_LOCK             : std_logic_vector(19 downto 0) := x"02300";
  constant REG_I2C_WR                         : std_logic_vector(19 downto 0) := x"02310";
  constant REG_I2C_RD                         : std_logic_vector(19 downto 0) := x"02320";
  constant REG_FPGA_CORE_TEMP                 : std_logic_vector(19 downto 0) := x"02330";
  constant REG_FPGA_CORE_VCCINT               : std_logic_vector(19 downto 0) := x"02340";
  constant REG_FPGA_CORE_VCCAUX               : std_logic_vector(19 downto 0) := x"02350";
  constant REG_FPGA_CORE_VCCBRAM              : std_logic_vector(19 downto 0) := x"02360";
  constant REG_FPGA_DNA                       : std_logic_vector(19 downto 0) := x"02370";
  constant REG_INT_TEST_4                     : std_logic_vector(19 downto 0) := x"02800";
  constant REG_INT_TEST_5                     : std_logic_vector(19 downto 0) := x"02810";

  --** Wishbone
  constant REG_WISHBONE_CONTROL               : std_logic_vector(19 downto 0) := x"04000";
  constant REG_WISHBONE_WRITE                 : std_logic_vector(19 downto 0) := x"04010";
  constant REG_WISHBONE_READ                  : std_logic_vector(19 downto 0) := x"04020";
  constant REG_WISHBONE_STATUS                : std_logic_vector(19 downto 0) := x"04030";
  -----------------------------------
  ---- GENERATED code END #1 ##  ----
  -----------------------------------

  --!
  --! --> CONTROL: Read/Write User Application Registers (Written by PCIe)
  ------------------------------------
  ---- ## GENERATED code BEGIN #2 ----
  ------------------------------------
  -- Bitfields of Control Record
  type bitfield_i2c_wr_t_type is record
    I2C_WREN                       : std_logic_vector(64 downto 64);  -- Any write to this register triggers an I2C read or write sequence
    WRITE_2BYTES                   : std_logic_vector(24 downto 24);  -- Write two bytes
    DATA_BYTE2                     : std_logic_vector(23 downto 16);  -- Data byte 2
    DATA_BYTE1                     : std_logic_vector(15 downto 8);   -- Data byte 1
    SLAVE_ADDRESS                  : std_logic_vector(7 downto 1);    -- Slave address
    READ_NOT_WRITE                 : std_logic_vector(0 downto 0);    -- READ/<o>WRITE</o>
  end record;

  type bitfield_i2c_rd_t_type is record
    I2C_RDEN                       : std_logic_vector(64 downto 64);  -- Any write to this register pops the last I2C data from the FIFO
  end record;

  type bitfield_wishbone_control_w_type is record
    WRITE_NOT_READ                 : std_logic_vector(32 downto 32);  -- wishbone write command wishbone read command
    ADDRESS                        : std_logic_vector(31 downto 0);   -- Slave address for Wishbone bus
  end record;

  type bitfield_wishbone_write_t_type is record
    WRITE_ENABLE                   : std_logic_vector(64 downto 64);  -- Any write to this register triggers a write to the Wupper to Wishbone fifo
    DATA                           : std_logic_vector(31 downto 0);   -- Wishbone
  end record;

  type bitfield_wishbone_read_t_type is record
    READ_ENABLE                    : std_logic_vector(64 downto 64);  -- Any write to this register triggers a read from the Wishbone to Wupper fifo
  end record;


  -- Control Record
  type register_map_control_type is record
    STATUS_LEDS                    : std_logic_vector(7 downto 0);    -- Board GPIO Leds
    LFSR_SEED_0                    : std_logic_vector(63 downto 0);   -- Least significant 64 bits of the LFSR seed
    LFSR_SEED_1                    : std_logic_vector(63 downto 0);   -- Bits 127 downto 64 of the LFSR seed
    LFSR_SEED_2                    : std_logic_vector(63 downto 0);   -- Bits 191 downto 128 of the LFSR seed
    LFSR_SEED_3                    : std_logic_vector(63 downto 0);   -- Bits 255 downto 192 of the LFSR seed
    APP_MUX                        : std_logic_vector(0 downto 0);    -- Switch between multiplier or LFSR.
                                                                      --   * 0 LFSR
                                                                      --   * 1 Loopback
                                                                      
    LFSR_LOAD_SEED                 : std_logic_vector(64 downto 64);  -- Writing any value to this register triggers the LFSR module to reset to the LFSR_SEED value
    APP_ENABLE                     : std_logic_vector(0 downto 0);    -- 1 Enables LFSR module or Loopback (depending on APP_MUX)
                                                                      -- 0 disable application
                                                                      
    I2C_WR                         : bitfield_i2c_wr_t_type;       
    I2C_RD                         : bitfield_i2c_rd_t_type;       
    INT_TEST_4                     : std_logic_vector(64 downto 64);  -- Fire a test MSIx interrupt #4
    INT_TEST_5                     : std_logic_vector(64 downto 64);  -- Fire a test MSIx interrupt #5
    WISHBONE_CONTROL               : bitfield_wishbone_control_w_type;
    WISHBONE_WRITE                 : bitfield_wishbone_write_t_type;
    WISHBONE_READ                  : bitfield_wishbone_read_t_type;
  end record;
  -----------------------------------
  ---- GENERATED code END #2 ##  ----
  -----------------------------------


  --!
  --! --> Read/Write User Application Registers DEFAULT values (Written by PCIe)
  ------------------------------------
  ---- ## GENERATED code BEGIN #3 ----
  ------------------------------------
  constant REG_STATUS_LEDS_C                       : std_logic_vector(7 downto 0)     := x"ab";                 -- Board GPIO Leds
  constant REG_LFSR_SEED_0_C                       : std_logic_vector(63 downto 0)    := x"0000000000000000";   -- Least significant 64 bits of the LFSR seed
  constant REG_LFSR_SEED_1_C                       : std_logic_vector(63 downto 0)    := x"0000000000000000";   -- Bits 127 downto 64 of the LFSR seed
  constant REG_LFSR_SEED_2_C                       : std_logic_vector(63 downto 0)    := x"0000000000000000";   -- Bits 191 downto 128 of the LFSR seed
  constant REG_LFSR_SEED_3_C                       : std_logic_vector(63 downto 0)    := x"0000000000000000";   -- Bits 255 downto 192 of the LFSR seed
  constant REG_APP_MUX_C                           : std_logic_vector(0 downto 0)     := "0";                   -- Switch between multiplier or LFSR.
                                                                                                                --   * 0 LFSR
                                                                                                                --   * 1 Loopback
                                                                                                                
  constant REG_LFSR_LOAD_SEED_C                    : std_logic_vector(64 downto 64)   := "0";                   -- Writing any value to this register triggers the LFSR module to reset to the LFSR_SEED value
  constant REG_APP_ENABLE_C                        : std_logic_vector(0 downto 0)     := "0";                   -- 1 Enables LFSR module or Loopback (depending on APP_MUX)
                                                                                                                -- 0 disable application
                                                                                                                
  constant REG_I2C_WR_I2C_WREN_C                   : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register triggers an I2C read or write sequence
  constant REG_I2C_WR_WRITE_2BYTES_C               : std_logic_vector(24 downto 24)   := "0";                   -- Write two bytes
  constant REG_I2C_WR_DATA_BYTE2_C                 : std_logic_vector(23 downto 16)   := x"00";                 -- Data byte 2
  constant REG_I2C_WR_DATA_BYTE1_C                 : std_logic_vector(15 downto 8)    := x"00";                 -- Data byte 1
  constant REG_I2C_WR_SLAVE_ADDRESS_C              : std_logic_vector(7 downto 1)     := "0000000";             -- Slave address
  constant REG_I2C_WR_READ_NOT_WRITE_C             : std_logic_vector(0 downto 0)     := "0";                   -- READ/<o>WRITE</o>
  constant REG_I2C_RD_I2C_RDEN_C                   : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register pops the last I2C data from the FIFO
  constant REG_INT_TEST_4_C                        : std_logic_vector(64 downto 64)   := "0";                   -- Fire a test MSIx interrupt #4
  constant REG_INT_TEST_5_C                        : std_logic_vector(64 downto 64)   := "0";                   -- Fire a test MSIx interrupt #5
  constant REG_WISHBONE_CONTROL_WRITE_NOT_READ_C   : std_logic_vector(32 downto 32)   := "0";                   -- wishbone write command wishbone read command
  constant REG_WISHBONE_CONTROL_ADDRESS_C          : std_logic_vector(31 downto 0)    := x"00000000";           -- Slave address for Wishbone bus
  constant REG_WISHBONE_WRITE_WRITE_ENABLE_C       : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register triggers a write to the Wupper to Wishbone fifo
  constant REG_WISHBONE_WRITE_DATA_C               : std_logic_vector(31 downto 0)    := x"00000000";           -- Wishbone
  constant REG_WISHBONE_READ_READ_ENABLE_C         : std_logic_vector(64 downto 64)   := "0";                   -- Any write to this register triggers a read from the Wishbone to Wupper fifo
  -----------------------------------
  ---- GENERATED code END #3 ##  ----
  -----------------------------------

  --!
  --! --> MONITOR: Read Only User Application Registers (Read by PCIe)
  ------------------------------------
  ---- ## GENERATED code BEGIN #4 ----
  ------------------------------------

--
-- GenericBoardInformation
--
  -- Bitfields of GenericBoardInformation
  type bitfield_generic_constants_r_type is record
    INTERRUPTS                     : std_logic_vector(15 downto 8);   -- Number of Interrupts
    DESCRIPTORS                    : std_logic_vector(7 downto 0);    -- Number of Descriptors
  end record;


  -- GenericBoardInformation
  type register_map_gen_board_info_type is record
    REG_MAP_VERSION                : std_logic_vector(15 downto 0);   -- Register Map Version, 1.0 formatted as 0x0100
    BOARD_ID_TIMESTAMP             : std_logic_vector(39 downto 0);   -- Board ID Date / Time in BCD format YYMMDDhhmm
    BOARD_ID_SVN                   : std_logic_vector(15 downto 0);   -- Board ID SVN Revision
    GENERIC_CONSTANTS              : bitfield_generic_constants_r_type;
    CARD_TYPE                      : std_logic_vector(63 downto 0);   -- Card Type:
                                                                      --   * 709 (0x2c5) VC709
                                                                      --   * 710 (0x2c6) HTG710
                                                                      --   * 711 (0x2c7) BNL711
                                                                      
end record;
--
-- HouseKeepingControlsAndMonitors
--
  -- Bitfields of HouseKeepingControlsAndMonitors
  type bitfield_i2c_wr_r_type is record
    I2C_FULL                       : std_logic_vector(25 downto 25);  -- I2C FIFO full
  end record;

  type bitfield_i2c_rd_r_type is record
    I2C_EMPTY                      : std_logic_vector(8 downto 8);    -- I2C FIFO Empty
    I2C_DOUT                       : std_logic_vector(7 downto 0);    -- I2C READ Data
  end record;


  -- HouseKeepingControlsAndMonitors
  type register_map_hk_monitor_type is record
    MMCM_MAIN_PLL_LOCK             : std_logic_vector(0 downto 0);    -- Main MMCM PLL Lock Status
    I2C_WR                         : bitfield_i2c_wr_r_type;       
    I2C_RD                         : bitfield_i2c_rd_r_type;       
    FPGA_CORE_TEMP                 : std_logic_vector(11 downto 0);   -- XADC temperature monitor for the FPGA CORE
                                                                      -- for Virtex7
                                                                      -- temp (C)= ((FPGA_CORE_TEMP* 503.975)/4096)-273.15
                                                                      -- for Kintex Ultrascale
                                                                      -- temp (C)= ((FPGA_CORE_TEMP* 502.9098)/4096)-273.8195
                                                                      
    FPGA_CORE_VCCINT               : std_logic_vector(11 downto 0);   -- XADC voltage measurement VCCINT = (FPGA_CORE_VCCINT *3.0)/4096
    FPGA_CORE_VCCAUX               : std_logic_vector(11 downto 0);   -- XADC voltage measurement VCCAUX = (FPGA_CORE_VCCAUX *3.0)/4096
    FPGA_CORE_VCCBRAM              : std_logic_vector(11 downto 0);   -- XADC voltage measurement VCCBRAM = (FPGA_CORE_VCCBRAM *3.0)/4096
    FPGA_DNA                       : std_logic_vector(63 downto 0);   -- Unique identifier of the FPGA
end record;
--
-- Wishbone
--
  -- Bitfields of Wishbone
  type bitfield_wishbone_write_r_type is record
    FULL                           : std_logic_vector(32 downto 32);  -- Wishbone
  end record;

  type bitfield_wishbone_read_r_type is record
    EMPTY                          : std_logic_vector(32 downto 32);  -- Indicates that the Wishbone to Wupper fifo is empty
    DATA                           : std_logic_vector(31 downto 0);   -- Wishbone read data
  end record;

  type bitfield_wishbone_status_r_type is record
    INT                            : std_logic_vector(4 downto 4);    -- interrupt
    RETRY                          : std_logic_vector(3 downto 3);    -- Interface is not ready to accept data cycle should be retried
    STALL                          : std_logic_vector(2 downto 2);    -- When pipelined mode slave can't accept additional transactions in its queue
    ACKNOWLEDGE                    : std_logic_vector(1 downto 1);    -- Indicates the termination of a normal bus cycle
    ERROR                          : std_logic_vector(0 downto 0);    -- Address not mapped by the crossbar
  end record;


  -- Wishbone
  type wishbone_monitor_type is record
    WISHBONE_WRITE                 : bitfield_wishbone_write_r_type;
    WISHBONE_READ                  : bitfield_wishbone_read_r_type;
    WISHBONE_STATUS                : bitfield_wishbone_status_r_type;
end record;
  

  -- Monitor interface toward the dma_control block
  type register_map_monitor_type is record
    register_map_gen_board_info  : register_map_gen_board_info_type;
    register_map_hk_monitor  : register_map_hk_monitor_type;
    wishbone_monitor  : wishbone_monitor_type;
  end record;
  -----------------------------------
  ---- GENERATED code END #4 ##  ----
  -----------------------------------

end package pcie_package ;

package body pcie_package is
    function to_sl( A: std_logic_vector) return std_logic is
    begin
        return A(A'low);
    end function to_sl;
end pcie_package;